library ieee;
use ieee.std_logic_1164.all;

entity regor is
port(
	ain, bin:in std_logic_vector(7 downto 0);
	sout:out std_logic_vector(7 downto 0)
);
end regor;

architecture dataflow of regor is
begin
	sout(0)<=(ain(0) or bin(0));
	sout(1)<=(ain(1) or bin(1));
	sout(2)<=(ain(2) or bin(2));
	sout(3)<=(ain(3) or bin(3));
	sout(4)<=(ain(4) or bin(4));
	sout(5)<=(ain(5) or bin(5));
	sout(6)<=(ain(6) or bin(6));
	sout(7)<=(ain(7) or bin(7));
end dataflow;